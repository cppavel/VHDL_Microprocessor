library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity control_memory is
    Port (FL : out std_logic; -- 0
            RZ : out std_logic; -- 1
            RN : out std_logic; -- 2
            RC : out std_logic; -- 3
            RV : out std_logic; -- 4
            MW : out std_logic; -- 5
            MM : out std_logic; -- 6
            RW : out std_logic; -- 7
            MD : out std_logic; -- 8
            FS : out std_logic_vector(4 downto 0); -- 9 to 13
            MB : out std_logic; -- 14
            TB : out std_logic; -- 15
            TA : out std_logic; -- 16
            TD : out std_logic; -- 17
            PL : out std_logic; -- 18
            PI : out std_logic; -- 19
            IL : out std_logic; -- 20
            MC : out std_logic; -- 21
            MS : out std_logic_vector(2 downto 0); -- 22 to 24
            NA : out std_logic_vector(16 downto 0); -- 25 to 41
            IN_CAR : in unsigned(16 downto 0));
end control_memory;

architecture Behavioral of control_memory is
    type mem_array is array(0 to 255) of std_logic_vector(41 downto 0);
    begin
    memory_m: process(IN_CAR)
    variable control_mem : mem_array:=(

-- | Next Address | MS    |M|I|P|P|T|T|T|M|     FS   |M|R|M|M|R|R|R|R|F|
-- | Next Address | MS    |C|L|I|L|D|A|B|B|     FS  |D|W|M|W|V|C|N|Z|L|
  
"000000000000000010010110000000000001000000",-- 0 IF 
"000000000111111110011000000000000000000000",-- 1 EX0 
"000000000000000000010000000100010010000001",-- 2 ADI 
"000000000000000000010000000000000110000000",-- 3 LD   
"000000000000000000010000000100001010000001",-- 4 INC
"000000000000000000010000000101110010000001",-- 5 NOT
"000000000000000000010000000000010010000001",-- 6 ADD
"000000000000000000010001000000000000000000",-- 7 BR
"000000000000010010010000000000000000000001",-- 8 BRZ (R[srcA] == 0, then branch)(8-10) Push value from reg through functional unit, get the flags
"000000000000001111000000000000000000000000",-- 9 - Go to BR if Z =1, else go to address a
"000000000000000000010000000000000000000000",-- a - Regardless go to IF
"000000000000011000010000100110000010000000",--  b - SR  Load the number of shifts into temp reg
"000000000000011010010000010000000000000001",--  c - Push the value through functional unit to get flags
"000000000000000001000000000000000000000000",--  d - if Z = 1 , go back to IF, otherwise increment
"000000000000011110010000000010100010000000",--  e - Shift right once 
"000000000000011010010000110000110010000001",--  f - decrement temp reg, go to state d to check the flag
    
    "000000000000000000000000000000000000000000",--  10
    "000000000000000000000000000000000000000000",--  11
    "000000000000000000000000000000000000000000",--  12
    "000000000000000000000000000000000000000000",--  13
    "000000000000000000000000000000000000000000",--  14
    "000000000000000000000000000000000000000000",--  15
    "000000000000000000000000000000000000000000",--  16
    "000000000000000000000000000000000000000000",--  17
    
    "000000000000000000000000000000000000000000",--  18
    "000000000000000000000000000000000000000000",--  19
    "000000000000000000000000000000000000000000",--  1a
    "000000000000000000000000000000000000000000",--  1b
    "000000000000000000000000000000000000000000",--  1c
    "000000000000000000000000000000000000000000",--  1d
    "000000000000000000000000000000000000000000",--  1e
    "000000000000000000000000000000000000000000",--  1f
    
    "000000000000000000000000000000000000000000",--  20
    "000000000000000000000000000000000000000000",--  21
    "000000000000000000000000000000000000000000",--  22
    "000000000000000000000000000000000000000000",--  23
    "000000000000000000000000000000000000000000",--  24
    "000000000000000000000000000000000000000000",--  25
    "000000000000000000000000000000000000000000",--  26
    "000000000000000000000000000000000000000000",--  27
    
    "000000000000000000000000000000000000000000",--  28
    "000000000000000000000000000000000000000000",--  29
    "000000000000000000000000000000000000000000",--  2a
    "000000000000000000000000000000000000000000",--  2b
    "000000000000000000000000000000000000000000",--  2c
    "000000000000000000000000000000000000000000",--  2d
    "000000000000000000000000000000000000000000",--  2e
    "000000000000000000000000000000000000000000",--  2f
    
    "000000000000000000000000000000000000000000",--  30
    "000000000000000000000000000000000000000000",--  31
    "000000000000000000000000000000000000000000",--  32
    "000000000000000000000000000000000000000000",--  33
    "000000000000000000000000000000000000000000",--  34
    "000000000000000000000000000000000000000000",--  35
    "000000000000000000000000000000000000000000",--  36
    "000000000000000000000000000000000000000000",--  37
    
    "000000000000000000000000000000000000000000",--  38
    "000000000000000000000000000000000000000000",--  39
    "000000000000000000000000000000000000000000",--  3a
    "000000000000000000000000000000000000000000",--  3b
    "000000000000000000000000000000000000000000",--  3c
    "000000000000000000000000000000000000000000",--  3d
    "000000000000000000000000000000000000000000",--  3e
    "000000000000000000000000000000000000000000",--  3f
    
    "000000000000000000000000000000000000000000",--  40
    "000000000000000000000000000000000000000000",--  41
    "000000000000000000000000000000000000000000",--  42
    "000000000000000000000000000000000000000000",--  43
    "000000000000000000000000000000000000000000",--  44
    "000000000000000000000000000000000000000000",--  45
    "000000000000000000000000000000000000000000",--  46
    "000000000000000000000000000000000000000000",--  47
    
    "000000000000000000000000000000000000000000",--  48
    "000000000000000000000000000000000000000000",--  49
    "000000000000000000000000000000000000000000",--  4a
    "000000000000000000000000000000000000000000",--  4b
    "000000000000000000000000000000000000000000",--  4c
    "000000000000000000000000000000000000000000",--  4d
    "000000000000000000000000000000000000000000",--  4e
    "000000000000000000000000000000000000000000",--  4f
    
    "000000000000000000000000000000000000000000",--  50
    "000000000000000000000000000000000000000000",--  51
    "000000000000000000000000000000000000000000",--  52
    "000000000000000000000000000000000000000000",--  53
    "000000000000000000000000000000000000000000",--  54
    "000000000000000000000000000000000000000000",--  55
    "000000000000000000000000000000000000000000",--  56
    "000000000000000000000000000000000000000000",--  57
    
    "000000000000000000000000000000000000000000",--  58
    "000000000000000000000000000000000000000000",--  59
    "000000000000000000000000000000000000000000",--  5a
    "000000000000000000000000000000000000000000",--  5b
    "000000000000000000000000000000000000000000",--  5c
    "000000000000000000000000000000000000000000",--  5d
    "000000000000000000000000000000000000000000",--  5e
    "000000000000000000000000000000000000000000",--  5f
    
    "000000000000000000000000000000000000000000",--  60
    "000000000000000000000000000000000000000000",--  61
    "000000000000000000000000000000000000000000",--  62
    "000000000000000000000000000000000000000000",--  63
    "000000000000000000000000000000000000000000",--  64
    "000000000000000000000000000000000000000000",--  65
    "000000000000000000000000000000000000000000",--  66
    "000000000000000000000000000000000000000000",--  67
    
    "000000000000000000000000000000000000000000",--  68
    "000000000000000000000000000000000000000000",--  69
    "000000000000000000000000000000000000000000",--  6a
    "000000000000000000000000000000000000000000",--  6b
    "000000000000000000000000000000000000000000",--  6c
    "000000000000000000000000000000000000000000",--  6d
    "000000000000000000000000000000000000000000",--  6e
    "000000000000000000000000000000000000000000",--  6f
    
    "000000000000000000000000000000000000000000",--  70
    "000000000000000000000000000000000000000000",--  71
    "000000000000000000000000000000000000000000",--  72
    "000000000000000000000000000000000000000000",--  73
    "000000000000000000000000000000000000000000",--  74
    "000000000000000000000000000000000000000000",--  75
    "000000000000000000000000000000000000000000",--  76
    "000000000000000000000000000000000000000000",--  77
    
    "000000000000000000000000000000000000000000",--  78
    "000000000000000000000000000000000000000000",--  79
    "000000000000000000000000000000000000000000",--  7a
    "000000000000000000000000000000000000000000",--  7b
    "000000000000000000000000000000000000000000",--  7c
    "000000000000000000000000000000000000000000",--  7d
    "000000000000000000000000000000000000000000",--  7e
    "000000000000000000000000000000000000000000",--  7f
    
    "000000000000000000000000000000000000000000",--  80
    "000000000000000000000000000000000000000000",--  81
    "000000000000000000000000000000000000000000",--  82
    "000000000000000000000000000000000000000000",--  83
    "000000000000000000000000000000000000000000",--  84
    "000000000000000000000000000000000000000000",--  85
    "000000000000000000000000000000000000000000",--  86
    "000000000000000000000000000000000000000000",--  87
    
    "000000000000000000000000000000000000000000",--  88
    "000000000000000000000000000000000000000000",--  89
    "000000000000000000000000000000000000000000",--  8a
    "000000000000000000000000000000000000000000",--  8b
    "000000000000000000000000000000000000000000",--  8c
    "000000000000000000000000000000000000000000",--  8d
    "000000000000000000000000000000000000000000",--  8e
    "000000000000000000000000000000000000000000",--  8f
    
    "000000000000000000000000000000000000000000",--  90
    "000000000000000000000000000000000000000000",--  91
    "000000000000000000000000000000000000000000",--  92
    "000000000000000000000000000000000000000000",--  93
    "000000000000000000000000000000000000000000",--  94
    "000000000000000000000000000000000000000000",--  95
    "000000000000000000000000000000000000000000",--  96
    "000000000000000000000000000000000000000000",--  97
    
    "000000000000000000000000000000000000000000",--  98
    "000000000000000000000000000000000000000000",--  99
    "000000000000000000000000000000000000000000",--  9a
    "000000000000000000000000000000000000000000",--  9b
    "000000000000000000000000000000000000000000",--  9c
    "000000000000000000000000000000000000000000",--  9d
    "000000000000000000000000000000000000000000",--  9e
    "000000000000000000000000000000000000000000",--  9f
    
    "000000000000000000000000000000000000000000",--  a0
    "000000000000000000000000000000000000000000",--  a1
    "000000000000000000000000000000000000000000",--  a2
    "000000000000000000000000000000000000000000",--  a3
    "000000000000000000000000000000000000000000",--  a4
    "000000000000000000000000000000000000000000",--  a5
    "000000000000000000000000000000000000000000",--  a6
    "000000000000000000000000000000000000000000",--  a7
    
    "000000000000000000000000000000000000000000",--  a8
    "000000000000000000000000000000000000000000",--  a9
    "000000000000000000000000000000000000000000",--  aa
    "000000000000000000000000000000000000000000",--  ab
    "000000000000000000000000000000000000000000",--  ac
    "000000000000000000000000000000000000000000",--  ad
    "000000000000000000000000000000000000000000",--  ae
    "000000000000000000000000000000000000000000",--  af
    
    "000000000000000000000000000000000000000000",--  b0
    "000000000000000000000000000000000000000000",--  b1
    "000000000000000000000000000000000000000000",--  b2
    "000000000000000000000000000000000000000000",--  b3
    "000000000000000000000000000000000000000000",--  b4
    "000000000000000000000000000000000000000000",--  b5
    "000000000000000000000000000000000000000000",--  b6
    "000000000000000000000000000000000000000000",--  b7
    
    "000000000000000000000000000000000000000000",--  b8
    "000000000000000000000000000000000000000000",--  b9
    "000000000000000000000000000000000000000000",--  ba
    "000000000000000000000000000000000000000000",--  bb
    "000000000000000000000000000000000000000000",--  bc
    "000000000000000000000000000000000000000000",--  bd
    "000000000000000000000000000000000000000000",--  be
    "000000000000000000000000000000000000000000",--  bf
    
    "000000000000000000000000000000000000000000",--  c0
    "000000000000000000000000000000000000000000",--  c1
    "000000000000000000000000000000000000000000",--  c2
    "000000000000000000000000000000000000000000",--  c3
    "000000000000000000000000000000000000000000",--  c4
    "000000000000000000000000000000000000000000",--  c5
    "000000000000000000000000000000000000000000",--  c6
    "000000000000000000000000000000000000000000",--  c7
    
    "000000000000000000000000000000000000000000",--  c8
    "000000000000000000000000000000000000000000",--  c9
    "000000000000000000000000000000000000000000",--  ca
    "000000000000000000000000000000000000000000",--  cb
    "000000000000000000000000000000000000000000",--  cc
    "000000000000000000000000000000000000000000",--  cd
    "000000000000000000000000000000000000000000",--  ce
    "000000000000000000000000000000000000000000",--  cf
    
    "000000000000000000000000000000000000000000",--  d0
    "000000000000000000000000000000000000000000",--  d1
    "000000000000000000000000000000000000000000",--  d2
    "000000000000000000000000000000000000000000",--  d3
    "000000000000000000000000000000000000000000",--  d4
    "000000000000000000000000000000000000000000",--  d5
    "000000000000000000000000000000000000000000",--  d6
    "000000000000000000000000000000000000000000",--  d7
    
    "000000000000000000000000000000000000000000",--  d8
    "000000000000000000000000000000000000000000",--  d9
    "000000000000000000000000000000000000000000",--  da
    "000000000000000000000000000000000000000000",--  db
    "000000000000000000000000000000000000000000",--  dc
    "000000000000000000000000000000000000000000",--  dd
    "000000000000000000000000000000000000000000",--  de
    "000000000000000000000000000000000000000000",--  df
    
    "000000000000000000000000000000000000000000",--  e0
    "000000000000000000000000000000000000000000",--  e1
    "000000000000000000000000000000000000000000",--  e2
    "000000000000000000000000000000000000000000",--  e3
    "000000000000000000000000000000000000000000",--  e4
    "000000000000000000000000000000000000000000",--  e5
    "000000000000000000000000000000000000000000",--  e6
    "000000000000000000000000000000000000000000",--  e7
    
    "000000000000000000000000000000000000000000",--  e8
    "000000000000000000000000000000000000000000",--  e9
    "000000000000000000000000000000000000000000",--  ea
    "000000000000000000000000000000000000000000",--  eb
    "000000000000000000000000000000000000000000",--  ec
    "000000000000000000000000000000000000000000",--  ed
    "000000000000000000000000000000000000000000",--  ee
    "000000000000000000000000000000000000000000",--  ef
    
    "000000000000000000000000000000000000000000",--  f0
    "000000000000000000000000000000000000000000",--  f1
    "000000000000000000000000000000000000000000",--  f2
    "000000000000000000000000000000000000000000",--  f3
    "000000000000000000000000000000000000000000",--  f4
    "000000000000000000000000000000000000000000",--  f5
    "000000000000000000000000000000000000000000",--  f6
    "000000000000000000000000000000000000000000",--  f7
    
    "000000000000000000000000000000000000000000",--  f8
    "000000000000000000000000000000000000000000",--  f9
    "000000000000000000000000000000000000000000",--  fa
    "000000000000000000000000000000000000000000",--  fb
    "000000000000000000000000000000000000000000",--  fc
    "000000000000000000000000000000000000000000",--  fd
    "000000000000000000000000000000000000000000",--  fe
    "000000000000000000000000000000000000000000");--  ff
        
        variable addr : integer;
        variable control_out : std_logic_vector(41 downto 0);
        
        begin
            addr := conv_integer(IN_CAR(7 downto 0));
            control_out := control_mem(addr);
            FL <= control_out(0) after 5 ns;
            RZ <= control_out(1) after 5 ns;
            RN <= control_out(2) after 5 ns;
            RC <= control_out(3) after 5 ns;
            RV <= control_out(4) after 5 ns;
            MW <= control_out(5) after 5 ns;
            MM <= control_out(6) after 5 ns;
            RW <= control_out(7) after 5 ns;
            MD <= control_out(8) after 5 ns;
            FS <= control_out(13 downto 9) after 5 ns;
            MB <= control_out(14) after 5 ns;
            TB <= control_out(15) after 5 ns;
            TA <= control_out(16) after 5 ns;
            TD <= control_out(17) after 5 ns;
            PL <= control_out(18) after 5 ns;
            PI <= control_out(19) after 5 ns;
            IL <= control_out(20) after 5 ns;
            MC <= control_out(21) after 5 ns;
            MS <= control_out(24 downto 22) after 5 ns;
            NA <= control_out(41 downto 25) after 5 ns;
        end process;
end Behavioral;


