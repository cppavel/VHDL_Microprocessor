library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity memory is 
    Port(address: unsigned(31 downto 0);
            write_data : in std_logic_vector(31 downto 0);
            MemWrite,Clk: in std_logic;
            read_data : out std_logic_vector(31 downto 0));
end memory;

architecture Behavioral of memory is

type mem_array is array(0 to 511) of std_logic_vector(31 downto 0);

begin
    mem_process: process (address, write_data, clk)
    variable data_mem : mem_array := (
    "00000000000000010000001000011111", "00000000000000011111110000000001",
    "00000000000000010000111111111111","00000000000000100000110001100000",
    "00000000000000101000110001100000","00000000000000110111111111100011",
    "00000000000000111000000000000010",X"00000000",
    X"00000000", "00000000000001000111111111110110", 
    "00000000000001011000110000000011","00000000000001000111110101010100",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"22891488",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000",
    X"00000000", X"00000000", X"00000000",X"00000000");
    variable addr:integer:=0;

    begin 
    if rising_edge(Clk)then
        addr:=conv_integer(unsigned(address(8 downto 0)));
        if MemWrite ='1' then
            data_mem(addr):=  write_data ;
        end if;
    end if;
    if MemWrite='0' then
         addr:=conv_integer(unsigned(address(8 downto 0)));
         read_data <= data_mem(addr) after 5 ns;
    end if;
    end process;
end Behavioral;
